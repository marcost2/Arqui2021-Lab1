module imem 
#(parameter N = 32) // name and default value
				(input logic [6:0] addr,
				 output logic [N-1:0] q);
		logic [N-1:0] ROM [128];

		initial 
           begin
           ROM = '{default:32'h00000000};
		     ROM [0:119] ='{32'hf8000286,
32'h8b1f03ff,
32'hab000000,
32'hf840028f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h54000100,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb4000dbf,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf800000f,
32'hab080000,
32'h54000101,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb4000c7f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf8000000,
32'h8b080000,
32'hab1e03de,
32'h54000102,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h54ffff63,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf800001e,
32'heb0103de,
32'h8b080000,
32'h54000104,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb40009bf,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf8000000,
32'hab080000,
32'h54000105,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb400087f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf8000000,
32'h8b080000,
32'hab1e03de,
32'h54000106,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h54ffff67,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf800001e,
32'h8b080000,
32'hab1e03de,
32'h54000108,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h54ffff69,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf800001e,
32'hab010021,
32'h5400010a,
32'h8b080000,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb400047f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf8000000,
32'heb030021,
32'h5400010b,
32'h8b080000,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb400033f,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf8000000,
32'hab020021,
32'h5400010c,
32'h8b080000,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb40001ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf8000000,
32'heb030063,
32'h5400010d,
32'h8b080000,
32'h8b1f03ff,
32'h8b1f03ff,
32'hb40000bf,
32'h8b1f03ff,
32'h8b1f03ff,
32'h8b1f03ff,
32'hf8000000,
32'hb400001f};







			  end
		always_comb
			begin
				q = ROM[addr];
			end
endmodule